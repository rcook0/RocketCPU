module boom_core_stub #(parameter int CORE_ID=0) (
  input  logic clk,
  input  logic reset_n
);
  // Placeholder for generated BOOM tile.
endmodule
